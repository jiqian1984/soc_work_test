`define DW 4
`define SP_Mult 4 
`define ONE_FRAME_LENGTH 1024